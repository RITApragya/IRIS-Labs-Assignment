/*
initial begin
	a = #5 2’d5;
	b = #5 2’d5;
	c = #5 2’d5;
*/

/*
initial begin
	a <= #5 2’d5;
	b <= #5 2’d5;
	c <= #5 2’d5;

*/


/*
a=1;b=2;c=3;
always @ (*) begin
	a = 5;
	b = a;
	c = a;
end 

*/


/*
a=1;b=2;c=3;
always @ (*) begin
	a <= 5;
	b <= a;
	c <= b;
end 

*/
